-- Pixel

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY majority_vote_circuit IS 
	PORT
	(
		B :  IN  STD_LOGIC;
		A :  IN  STD_LOGIC;
		C :  IN  STD_LOGIC;
		Y :  OUT  STD_LOGIC;
	);
END majority_vote_circuit;

ARCHITECTURE bdf_type OF majority_vote_circuit IS 

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;


BEGIN 



SYNTHESIZED_WIRE_0 <= A AND B;


SYNTHESIZED_WIRE_1 <= A AND C;


SYNTHESIZED_WIRE_2 <= C AND B;


SYNTHESIZED_WIRE_3 <= SYNTHESIZED_WIRE_0 XOR SYNTHESIZED_WIRE_1;


Y <= SYNTHESIZED_WIRE_3 XOR SYNTHESIZED_WIRE_2

END bdf_type;